//A 4-core system!
`define NUM_CORES 4
`define CORE_IDX_WIDTH 2
